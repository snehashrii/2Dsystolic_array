(*synthesize*)
module trial(Empty);

Reg#(int) cyc <- mkReg(0);

rule kjhjh;

cyc<=3000;
$display("%0d", cyc);

endrule

endmodule